library ieee;
use ieee.std_logic_1164.all;
use work.inv_MixColumns_package.all;
use work.inv_ShiftRows_package.all;
use work.inv_SubBytes_package.all;

entity MixColumns_tb is
end MixColumns_tb;

architecture arch of MixColumns_tb is
   
   
   signal input, output : std_logic_vector (127 downto 0);
   
begin

  input <= inv_MixColumns(x"5f72641557f5bc92f7be3b291db9f91a");
  
end arch ; 